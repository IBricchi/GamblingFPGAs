module Testing (
input in,
output out
);

reg internal = 1;

assign out = in;

endmodule